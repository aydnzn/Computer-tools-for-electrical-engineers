** Profile: "SCHEMATIC1-circuitwithopampsusingVCVS"  [ C:\USERS\AYD�N UZUN\circuitwithopampsusingvcvs-PSpiceFiles\SCHEMATIC1\circuitwithopampsusingVCVS.sim ] 

** Creating circuit file "circuitwithopampsusingVCVS.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "C:/Cadence/SPB_17.2/tools/capture/library/pspice/userlib/ad8608.lib" 
* From [PSPICE NETLIST] section of C:\Users\Ayd�n Uzun\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 10s 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
